//tb for route computation unit 
import params_noc::*;
module route_computation_tb()();

endmodule