
module status_Buffer #(parameter BUFFER_SIZE = 8)

();


endmodule