import params_noc::*;

//Status Buffer verilog code which tells us about the status of the current flit 
module status_Buffer #(parameter BUFFER_SIZE = 8)

(
  input clk,					                            //clk
  input rst_n,					                          //reset
  input read_i,					                          //read signal 
  input write_i,				                          //write signal
  output logic buf_empty,			                    //buffer empty
  output logic buf_full,			                    //buffer full
  output logic buf_On_Off,			                  //Buffer on and off signal 
  input flit_Data_noVC input_Data,	              //input flit without vc info
  output flit_Data_withvc output_Data,		        //output flit after being assigned to a vc 
  input inout_Port port_i,			                  //input port
  output inout_Port port_o,			                  //output port 
  input [VC_Size-1:0] vc_New,			                //Vc allocation 
  input vc_Val,					                          //Vc valid 
  output logic vc_Req,				                    //Vc allocationn request
  output logic vc_Alloc,			                    //Vc allocation for the next flit sent to the upstream router 
  output logic switch_Req,			                  // switch allocation request
  output logic err,				                        //error
  output logic [VC_Size-1:0] downstream_Vc	      //signal to tell if vc is available in down stream router 
);

  
  logic [VC_Size-1:0] downstream_Vc_Next;
  logic read_Cmd, write_Cmd;
  logic end_Packet, end_Packet_Next;
  logic vc_Alloc_next;
  logic err_Next;
  flit_Data_noVC read_flit;
  inout_Port port_o_Next;
  
  typedef enum logic [1:0]{IDLE, VC, SWITCH} state_t;
  state_t p_state, nxt_state;

always@(posedge clk, negedge rst_n) begin 
  if(!rst_n)begin
    p_state 		<= IDLE;
    port_o  		<= LOCAL;
    downstream_Vc     	<= 0;
    end_Packet          <= 0;
    vc_Alloc    	<= 0;
    err             	<= 0;
  end
  else begin
    p_state 		<= nxt_state;
    port_o          	<= port_o_Next;
    downstream_Vc     	<= downstream_Vc_Next;
    end_Packet          <= end_Packet_Next;
    vc_Alloc    	<= vc_Alloc_next;
    err             	<= err_Next;
  end
end 
    

//Circular Buffer instantiation
circular_Buffer #(.BUFFER_SIZE(BUFFER_SIZE)) cirbuf (.clk(clk), .rst_n(rst_n), .input_Data(input_Data), .output_Data(output_Data), .read_i(read_i), .write_i(write_i),
  .buf_empty(buf_empty), .buf_full(buf_full), .buf_On_Off(buf_On_Off));

// //FSM logic 
// always@(*) begin 

//   case(state_t)
//     default: begin 
//     end 
//     IDLE: begin 
//     end 
//     VC: begin 
//     end 
//     SWITCH: begin 
//     end 
//   endcase
// end

endmodule